// 
module ALU(srcA, srcB, ALUop, result, ALUzero);
input[31:0] srcA, srcB;
input ALUop;
output [31:0] result, ALUzero;


endmodule