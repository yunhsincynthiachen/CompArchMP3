module pc_we_handler(ALUzero_out, pc_we, handler_out);
input[31:0] ALUzero_out;
input pc_we;
output handler_out;

//oring the last bit of ALUzero_out with pc_we

endmodule  