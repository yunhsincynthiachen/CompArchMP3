module TwoInputMuxes(wordA, wordB, control_signal, output_twoinput);
input[31:0] wordA, wordB;
input control_signal;
output[31:0] output_twoinput;

endmodule 