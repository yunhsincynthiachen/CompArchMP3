module signextend(imm16_ir, signextend_out);
input[15:0] imm16_ir; 
output[15:0] signextend_out;

endmodule 