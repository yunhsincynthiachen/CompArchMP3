module Value4(four_out);
output[31:0] four_out;
assign four_out = 'b00000000000000000000000000000100;

endmodule 