module value31(register_out);
output[4:0] register_out = 'b11111;

endmodule 