module value4(four_out);
output[31:0] four_out = 0x04;

endmodule 